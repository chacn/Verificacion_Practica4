module Serial_equalizer{
	//Input ports.
	input clk,
	input reset,
	input LRC_signal,
	input left_data,
	input right_data,
	
	//Output ports.
	output

}


endmodule 